module uart_rx (
    input clk,
    input rst_n,
    input uart_rx,

    output [7:0] rx_data,
    output rx_valid
);

    // TODO: UART 接收实现

endmodule