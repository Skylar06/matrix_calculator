module led_status (
    input clk,
    input rst_n,
    input error_flag,
    input busy_flag,
    input done_flag,

    output [2:0] led
);

    // TODO: LED效果

endmodule