module matrix_top (
    input clk,
    input rst_n,
    input [7:0] sw,
    input [3:0] key,
    input uart_rx,

    output uart_tx,
    output [2:0] led,
    output [3:0] seg_sel,
    output [7:0] seg_data
);

    // TODO: 声明内部连线，并实例化下面 9 个子模块

endmodule