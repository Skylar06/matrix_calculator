module uart_tx (
    input clk,
    input rst_n,
    input tx_start,
    input [7:0] tx_data,

    output uart_tx
);

    // TODO: UART 发送实现

endmodule